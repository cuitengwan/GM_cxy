`timescale 1ns/1ns
module aaa();
    reg clk;
    reg rstn;
    reg[2047:0] din;
    reg start;
    wire[1023:0] dout;
    wire valid;
    sm3top sm3top(clk,rstn,din,start,dout,valid);
    always @* begin
        #5 clk <= ~clk;
    end
    initial begin
        clk <= 0;
        rstn <= 0;
        start <= 0;
        /*
        din[2047:1536] <= 512'h0;
        din[1535:1024] <= 512'hx;
        din[1023:512]  <= 512'h0;
        din[511:0]     <= 512'hz;
        */
        din <= 0;
        #20;
        rstn <= 1;
        #40;
        
        // din[2047:2016] <= 32'h61626380;
        // din[1567:1536] <= 32'h00000018;
        /*
        din[1535:1504] <= 32'h61626380;
        din[1055:1024] <= 32'h00000018;
        
        din[1023:992] <= 32'h61626380;
        din[543:512] <= 32'h00000018;
        din[511:480] <= 32'h61626380;
        din[31:0] <= 32'h00000018;
        */
        din[2047:1536] <= 512'h61626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364;

        din[1535:1024] <= 512'h61626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364;

        din[1023:512] <= 512'h61626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364;

        din[511:0] <= 512'h61626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364616263646162636461626364;

        
        start <= 1;
        #10;
        //din <= 0;
        start <= 0;

        #3500;
        din[2047:1536] <= 512'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200;
        din[1535:1024] <= 512'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200;
        din[1023:512] <= 512'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200;
        din[511:0] <= 512'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200;
        start <= 1;
        #10;
        start <= 0;

    end
endmodule
